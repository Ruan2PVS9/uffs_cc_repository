library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity batalhaNaval_ruan is
    port(
        SW: in std_logic_vector(9 downto 0);
        key: in std_logic_vector(3 downto 0);

        LEDG: out std_logic_vector(6 downto 0);
        LEDR: out std_logic_vector(9 downto 0);
        hex0: out std_logic_vector(6 downto 0);
        hex1: out std_logic_vector(6 downto 0);
        hex2: out std_logic_vector(6 downto 0);
        hex3: out std_logic_vector(6 downto 0)
        
    );
end batalhaNaval_ruan;

architecture main of batalhaNaval_ruan is

    type estado is (set, shot,win,lost);

    signal state : estado := set;

    -- variable cont_erros : std_logic_vector(2 downto 0) := "000";
    -- variable cont_acertos : std_logic_vector(1 downto 0) := "00";
    -- variable cont_disparos : std_logic_vector(3 downto 0) := "0000";
    -- -- '-' para representar um estado não inicializado.
    -- variable nav1, nav2_casa1, nav2_casa2 : std_logic_vector(3 downto 0) := "----";
    -- variable decod_disp, cod_disp : std_logic_vector(3 downto 0);


    function codificar(decodificado : std_logic_vector(3 downto 0)) return std_logic_vector is
        variable A, B, C, D : std_logic;
        variable resultado : std_logic_vector(3 downto 0);
    begin
        A := decodificado(3);
        B := decodificado(2);
        C := decodificado(1);
        D := decodificado(0);

        -- a = ~B⋅~C⋅~D + ~A⋅~B⋅C⋅D + ~A⋅B⋅~C⋅D + B⋅C⋅~D + A⋅~D
        resultado(3) := (   (not B and not C and not D) or
                            (not A and not B and C and D) or 
                            (not A and b and not C and D ) or 
                            (B and C and not D) or 
                            (A and not D)
                        );

        -- b = ~A⋅~B⋅D + ~A⋅C + ~B⋅C + C⋅~D
        resultado(2) := (   (not A and not B and D) or 
                            (not A and C) or 
                            (not B and C) or 
                            (c and not D) 
                        );
        
        -- c = ~A⋅~D + ~B⋅~D + A⋅C⋅D
        resultado(1) := (   (not A and not D) or 
                            (not B and not D) or 
                            (A and C and D) 
                        );

        -- d = ~A⋅~B⋅C + ~A⋅C⋅D + A⋅~B⋅~D + A⋅~C⋅~D + A⋅B⋅~C + B⋅C⋅D
        resultado(0) := (   (not A and not B and C) or 
                            (not A and C and D) or 
                            (A and not B and not D) or 
                            (A and not C and not D) or 
                            (A and B and not C) or 
                            (B and C and D) 
                        );

        return resultado;
    end codificar;

    function decodificar(codificado : std_logic_vector(3 downto 0)) return std_logic_vector is
        variable a, b, c, d : std_logic;
        variable resultado : std_logic_vector(3 downto 0);
    begin
        a := codificado(3);
        b := codificado(2);
        c := codificado(1);
        d := codificado(0);
        -- A = ~a⋅~b⋅~c + ~b⋅d + ~a⋅b⋅c⋅~d + a⋅b⋅~c⋅~d + a⋅c⋅d
        resultado(3) := (   (not a and not b and not c) or
                            (not b and d) or
                            (not a and b and c and not d) or
                            (a and b and not c and not d) or
                            (a and c and d) 
                        );

        -- B = ~a⋅~b⋅c + ~a⋅~c⋅d + a⋅~b⋅~c + a⋅b⋅~d
        resultado(2) := (   (not a and not b and c) or
                            (not a and not c and d) or
                            (a and not b and not c) or
                            (a and b and not d)
                        );

        -- C = ~a⋅c⋅d + b⋅d + b⋅c
        resultado(1) := (   (not a and c and d) or
                            (b and d) or
                            (b and c) 
                        );

        -- D = ~a⋅~b⋅d + ~b⋅~c⋅~d + ~a⋅b⋅~d + b⋅~c⋅d
        resultado(0) := (   (not a and not b and d) or
                            (not b and not c and not d) or
                            (not a and b and not d) or
                            (b and not c and d)
                        );

        return resultado;
    end decodificar;

    -- function set_casa2(cod_casa1 : std_logic_vector(3 downto 0); v_or_h : std_logic) return std_logic_vector is
    --     variable cod_casa2 : std_logic_vector(3 downto 0);
    --     variable decod_casa_1 : std_logic_vector(3 downto 0);
    --     variable decod_casa_2 : std_logic_vector(3 downto 0);
    -- begin
    --     decod_casa_1 := decodificar(cod_casa1);
    --     if (v_or_h = "0") then
    --         if decod_casa_1 = "0011" then
    --             decod_casa_2 := "0010";
    --         elsif decod_casa_1 = "0111" then
    --             decod_casa_2 := "0110";
    --         elsif decod_casa_1 = "1011" then
    --             decod_casa_2 := "1010";
    --         elsif decod_casa_1 = "1111" then
    --             decod_casa_2 := "1110";
    --         else
    --             decod_casa_2 := decod_casa_1 + "0001";
    --         end if ;
    --     elsif (v_or_h = "1") then
    --         if decod_casa_1 = "1100" then
    --             decod_casa_2 := "1000";
    --         elsif decod_casa_1 = "1101" then
    --             decod_casa_2 := "1001";
    --         elsif decod_casa_1 = "1110" then
    --             decod_casa_2 := "1010";
    --         elsif decod_casa_1 = "1111" then
    --             decod_casa_2 := "1011";
    --         else
    --             decod_casa_2 := decod_casa_1 + "0100";
    --         end if ;
    --     end if ;
    --     cod_casa2 := codificar(decod_casa_2);
    --     return cod_casa2;
    -- end set_casa2;
    
begin
    -- variable cont_erros : std_logic_vector(2 downto 0) := "000";
    -- variable cont_acertos : std_logic_vector(1 downto 0) := "00";
    -- variable cont_disparos : std_logic_vector(3 downto 0) := "0000";
    -- -- '-' para representar um estado não inicializado.
    -- variable nav1, nav2_casa1, nav2_casa2 : std_logic_vector(3 downto 0) := "----";
    -- variable decod_disp, cod_disp : std_logic_vector(3 downto 0);

    process(key(0), key(1))

    -- variable cont_erros : std_logic_vector(2 downto 0) := "000";
    -- variable cont_acertos : std_logic_vector(1 downto 0) := "00";
    -- variable cont_disparos : std_logic_vector(3 downto 0) := "0000";


    variable cont_erros : std_logic_vector(2 downto 0) := "000";
    variable cont_acertos : std_logic_vector(1 downto 0) := "00";
    variable cont_disparos : std_logic_vector(3 downto 0) := "0000";
    -- '-' para representar um estado não inicializado.
    variable nav1, nav2_casa1, nav2_casa2 : std_logic_vector(3 downto 0) := "----";
    variable decod_disp, cod_disp : std_logic_vector(3 downto 0);
    variable decod_casa_1, decod_casa_2 : std_logic_vector(3 downto 0) := "----";
    variable somar3 :std_logic_vector(3 downto 0) ;
    variable somar1 :std_logic_vector(1 downto 0) ;
    variable somar2 :std_logic_vector(2 downto 0) ;

    begin

    if (key(1) = '0') then
        
        cont_erros := "000";
        cont_acertos := "00";
        cont_disparos := "0000";

        nav1 := "----";
        nav2_casa1 := "----";
        nav2_casa2 := "----";

        ledg <= "1111111";
        ledr <= "1111111111";
        ledr <= "0000000000";
        ledg <= "0000000";


    elsif (key(0)'EVENT and key(0) = '0') then
        if (state = set) then
            if (sw(4) = '0' and key(2) = '0') then
                -- set1 = 
                -- hex <= "0123456"

                hex3 <= "1011011";
                hex2 <= "1001111";
                hex1 <= "0001111";
                hex0 <= "1001111";

                nav1(0) := sw(0);
                nav1(1) := sw(1);
                nav1(2) := sw(2);
                nav1(3) := sw(3);
                ledg(0) <= '1';
            elsif (sw(4) = '1' and key(2) = '0') then
                -- set2 = 
                -- hex <= "0123456"

                hex3 <= "1011011";
                hex2 <= "1001111";
                hex1 <= "0001111";
                hex0 <= "1101101";

                nav2_casa1(0) := sw(0);
                nav2_casa1(1) := sw(1);
                nav2_casa1(2) := sw(2);
                nav2_casa1(3) := sw(3);
                ledg(1) <= '1';


                decod_casa_1 := decodificar(nav2_casa1);
                if (sw(6) = '0') then
                    -- nav2_casa2 <= set_casa2(nav2_casa1,"0");
                    if (decod_casa_1 = "0011") then
                        decod_casa_2 := "0010";
                    elsif (decod_casa_1 = "0111") then
                        decod_casa_2 := "0110";
                    elsif (decod_casa_1 = "1011") then
                        decod_casa_2 := "1010";
                    elsif (decod_casa_1 = "1111") then
                        decod_casa_2 := "1110";
                    else
                        somar3 := "0001";
                        decod_casa_2 := std_logic_vector(unsigned(decod_casa_1) + unsigned(somar3));
                    end if ;
                elsif (sw(6) = '1') then
                    -- nav2_casa2 <= set_casa2(nav2_casa1,"1");
                    if (decod_casa_1 = "1100") then
                        decod_casa_2 := "1000";
                    elsif (decod_casa_1 = "1101") then
                        decod_casa_2 := "1001";
                    elsif (decod_casa_1 = "1110") then
                        decod_casa_2 := "1010";
                    elsif (decod_casa_1 = "1111") then
                        decod_casa_2 := "1011";
                    else
                        somar3 := "0100";
                        decod_casa_2 := std_logic_vector(unsigned(decod_casa_1) + unsigned(somar3));
                    end if ;
                end if;
                if (nav2_casa2 /= "----") then
                    nav2_casa2 := codificar(decod_casa_2);
                    ledg(2) <= '1';
                end if;
            end if;
            if ((nav1 /= "----") and (nav2_casa1 /= "----") and (nav2_casa2 /= "----") and (sw(5) = '1')) then
                state <= shot;
            end if ;
        elsif (state = shot) then
            decod_disp(0) := sw(0);
            decod_disp(1) := sw(1);
            decod_disp(2) := sw(2);
            decod_disp(3) := sw(3);
            if (key(2) = '0') then
                -- disX = 
                -- hex <= "0123456"

                hex3 <= "1111110";
                hex2 <= "1111001";
                hex1 <= "1011011";
                case cont_disparos is
                    when "0000" =>
                        hex0 <= "1001111";

                    when "0001" =>
                        hex0 <= "1101101";

                    when "0010" =>
                        hex0 <= "1101101";

                    when others =>
                        -- cont_erros <= cont_erros + "001";
                        ledr <= "1111111111";
                end case;
                -- hex0 <= "0123456";

                cod_disp := codificar(decod_disp);

                if (cod_disp = nav1) then
                    ledg(0) <= '0';
                    somar1 := "01";
                    cont_acertos := std_logic_vector(unsigned(cont_acertos) + unsigned(somar1));
                elsif (cod_disp = nav2_casa1) then
                    ledg(1) <= '0';
                    somar1 := "01";
                    cont_acertos := std_logic_vector(unsigned(cont_acertos) + unsigned(somar1));
                elsif (cod_disp = nav2_casa2) then
                    ledg(2) <= '0';
                    somar1 := "01";
                    cont_acertos := std_logic_vector(unsigned(cont_acertos) + unsigned(somar1));
                else
                    somar2 :="001";
                    cont_erros := std_logic_vector(unsigned(cont_erros) + unsigned(somar2));
                    
                end if ;
                somar3 := "0001";
                cont_disparos := std_logic_vector(unsigned(cont_disparos) + unsigned(somar2));
                
            end if;
            if (cont_acertos = "11") then
                state <= lost;
            
            elsif (cont_acertos = "110") then
                state <= win;
                
            end if ;
        end if;
    end if ;
    end process;
    process(state)
    begin
        if (state = win) then
            ledg <= "1111111";
            ledr <= "0000000000";
        elsif (state = lost) then
            ledg <= "0000000";
            ledr <= "1111111111";
            
        end if ;

    end process;



end architecture;